library verilog;
use verilog.vl_types.all;
entity counterDIv_vlg_vec_tst is
end counterDIv_vlg_vec_tst;
