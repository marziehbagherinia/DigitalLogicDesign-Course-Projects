library verilog;
use verilog.vl_types.all;
entity CounterDivider_vlg_vec_tst is
end CounterDivider_vlg_vec_tst;
