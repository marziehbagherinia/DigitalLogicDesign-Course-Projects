library verilog;
use verilog.vl_types.all;
entity CounterDivider_tst is
end CounterDivider_tst;
