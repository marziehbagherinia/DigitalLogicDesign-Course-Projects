library verilog;
use verilog.vl_types.all;
entity controllerTB is
end controllerTB;
