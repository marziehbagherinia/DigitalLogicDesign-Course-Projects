`timescale 1 ps/ 1 ps

module square_wave(clk,
                   rst,
                   counter,
                   square_out);
                   
   input clk,
         rst;
   input [7:0]  counter;
   output reg [7:0] square_out;

   always @(posedge clk) begin
        if (rst == 1'b0  &&  counter < 8'b10000000)
          square_out <= 8'b11111111;
        else
          square_out <= 8'b0;
   end

endmodule