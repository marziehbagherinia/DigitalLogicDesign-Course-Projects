library verilog;
use verilog.vl_types.all;
entity testTB is
end testTB;
