library verilog;
use verilog.vl_types.all;
entity CounterDivider_vlg_check_tst is
    port(
        cout            : in     vl_logic;
        MaxMin2         : in     vl_logic;
        out0            : in     vl_logic;
        out1            : in     vl_logic;
        out2            : in     vl_logic;
        out3            : in     vl_logic;
        out4            : in     vl_logic;
        out5            : in     vl_logic;
        out6            : in     vl_logic;
        out7            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end CounterDivider_vlg_check_tst;
