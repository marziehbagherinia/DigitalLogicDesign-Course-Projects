library verilog;
use verilog.vl_types.all;
entity CA5TB is
end CA5TB;
