library verilog;
use verilog.vl_types.all;
entity WaveformGenerator_vlg_vec_tst is
end WaveformGenerator_vlg_vec_tst;
